`include "counter.sv"
